module 2mux
	(
	// ------------------------------------------------------------ 
	// Inputs
	// ------------------------------------------------------------
	input [15:0] data,
	input select,
	// ------------------------------------------------------------

	// ------------------------------------------------------------ 
	// Outputs
	// ------------------------------------------------------------
	output [15:0] out
	// ------------------------------------------------------------ 
	);

// -------------------------------------------------------------------- 
// Logic Declaration
// --------------------------------------------------------------------	
	always @(*) begin
	
		out = data[select];

	end
// --------------------------------------------------------------------
endmodule
// --------------------------------------------------------------------

