module mux8
	(
	// ------------------------------------------------------------ 
	// Inputs
	// ------------------------------------------------------------
	input [15:0] data0,
	input [15:0] data1,
	input [15:0] data2,
	input [15:0] data3,
	input [15:0] data4,
	input [15:0] data5,
	input [15:0] data6,
	input [15:0] data7,
	input [2:0]select,
	// ------------------------------------------------------------

	// ------------------------------------------------------------ 
	// Outputs
	// ------------------------------------------------------------
	output [15:0] out
	// ------------------------------------------------------------ 
	);

// -------------------------------------------------------------------- 
// Logic Declaration
// --------------------------------------------------------------------	
	always @(*) begin

		case(select)
			3'b000: begin
				out = data0;
			end
			3'b001: begin
				out = data1;
			end
			3'b010: begin
				out = data2;
			end
			3'b011: begin
				out = data3;
			end
			3'b100: begin
				out = data4;
			end
			3'b101: begin
				out = data5;
			end
			3'b110: begin
				out = data6;
			end
			3'b111: begin
				out = data7;
			end
		endcase

	end
// --------------------------------------------------------------------
endmodule
// --------------------------------------------------------------------

