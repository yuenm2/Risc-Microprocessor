module pc (
	// ------------------------------------------------------------ 
	// Inputs
	// ------------------------------------------------------------
	input wire clk,
	input wire[15:0] pc_i,
	// ------------------------------------------------------------

	// ------------------------------------------------------------ 
	// Outputs
	// ------------------------------------------------------------
	output reg[15:0] pc_o
	// ------------------------------------------------------------ 
	);
	
	always @(posedge clk) begin
		pc_o <= pc_i;
	end

endmodule
// --------------------------------------------------------------------